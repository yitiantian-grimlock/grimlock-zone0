//test for vscode and github
